cdl/uart03.cdl