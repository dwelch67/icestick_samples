cdl/uart02.cdl