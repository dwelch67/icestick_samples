
module blinker01
(
    clock clk,
    output bit LED1,
    output bit LED2,
    output bit LED3,
    output bit LED4,
    output bit LED5,
    output bit RS232_Tx,
    input bit PMOD1,
    input bit PMOD2,
    input bit PMOD3,
    input bit PMOD4
)
{
    default clock clk;
    default reset active_high PMOD4 ;

    clocked bit[32] XCOUNT = 0;
    clocked bit[8] UCOUNT = 0;
    clocked bit[1] UARTTX = 0;

    the_code:
    {
        XCOUNT <= XCOUNT + 1;

        LED1 = XCOUNT[23];
        LED2 = XCOUNT[23];
        LED3 = XCOUNT[23];
        LED4 = XCOUNT[23];
        LED5 = XCOUNT[23];

        if(UCOUNT == 103)
        {
            UCOUNT <= 0;
            UARTTX <= UARTTX + 1;
        }
        else
        {
            UCOUNT <= UCOUNT + 1;
        }
        RS232_Tx = UARTTX;
    }
}
