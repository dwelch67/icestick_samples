
//cdl --model csram --cpp csram.cpp csram.cdl

extern module csram
(
    input   bit[1]  in_output_enable,
    input   bit[1]  in_write_enable,
    input   bit[16] in_address,
    input   bit[16] in_data,
    output  bit[16] out_data
)
{
    timing comb input in_output_enable;
    timing comb input in_write_enable;
    timing comb input in_address;
    timing comb input in_data;
    timing comb output out_data;
}

module csram
(
    input   bit[1]  in_output_enable,
    input   bit[1]  in_write_enable,
    input   bit[16] in_address,
    input   bit[16] in_data,
    output  bit[16] out_data
)
{
    sram_code:
    {
        out_data = 16hFFFF;
        if(in_output_enable==1b1)
        {
            full_switch(in_address)
            { //0001 0000 0100 0001
                //case 16h3000: { out_data = 0x9040; }
                //case 16h3001: { out_data = 0x5060; }
                //case 16h3002: { out_data = 0x1027; }
                //case 16h3003: { out_data = 0x103F; }
                //case 16h3004: { out_data = 0x0BFE; }
                //case 16h3005: { out_data = 0xF025; }
                //case 16h3006: { out_data = 0x0FF9; }
include "program.cdl"
                default: { out_data = 0xFFFF; }
            }
        }
        if(in_write_enable==1b1)
        {
            out_data = in_data;
        }
    }
}

