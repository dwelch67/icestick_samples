extern module csram
(
    input   bit[1]  in_output_enable,
    input   bit[1]  in_write_enable,
    input   bit[16] in_address,
    input   bit[16] in_data,
    output  bit[16] out_data
)
{
    timing comb input in_output_enable;
    timing comb input in_write_enable;
    timing comb input in_address;
    timing comb input in_data;
    timing comb output out_data;
}

extern module core
(
    clock          clock_in,
    input  bit     reset_in,

    input  bit[16] mem_in,
    output bit[16] mem_out,
    output bit[16] mem_add,
    output bit[1]  mem_oe,
    output bit[1]  mem_we,
    output bit[1]  mem_fetch,
    output bit[8]  led_out
)
{
    timing to rising clock clock_in reset_in;
    timing to rising clock clock_in mem_in;
    timing from rising clock clock_in mem_out;
    timing from rising clock clock_in mem_add;
    timing from rising clock clock_in mem_oe;
    timing from rising clock clock_in mem_we;
    timing from rising clock clock_in mem_fetch;
    timing from rising clock clock_in led_out;
}

module top
(
    clock          in_clock,
    input  bit     in_reset,
    output bit[8]   out_led
)
{
    default clock in_clock ;
    default reset active_high in_reset ;

    net  bit[8] net_led_out;
    net bit[1] net_mem_fetch;

    net bit net_output_enable;
    net bit net_write_enable;
    net bit[16] net_address;
    net bit[16] net_in_data;
    net bit[16] net_out_data;

    top_code:
    {
        csram mem
        (
            in_output_enable    <= net_output_enable,
            in_write_enable     <= net_write_enable,
            in_address          <= net_address,
            in_data             <= net_in_data,
            out_data            => net_out_data
        );
        core core0
        (
            clock_in <- in_clock,
            reset_in <= in_reset,

            mem_in <= net_out_data,
            mem_oe => net_output_enable,
            mem_we => net_write_enable,
            mem_add => net_address,
            mem_out => net_in_data,
            mem_fetch => net_mem_fetch,
            led_out => net_led_out
        );
        out_led = net_led_out;
    }
}
