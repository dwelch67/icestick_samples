
module blinker02
(
    clock clk,
    output bit LED0,
    output bit LED1,
    output bit LED2,
    output bit LED3,
    output bit LED4,
    output bit LED5,
    output bit LED6,
    output bit LED7,
    input bit NOTRESET
)
{
    default clock clk;
    default reset active_high NOTRESET ;
    clocked bit[12] XCOUNT = 1;
    clocked bit[12] ZCOUNT = 0x10;
    clocked bit ledout = 0;
    clocked bit state = 0;
    
    the_code:
    {
        XCOUNT <= XCOUNT + 1;

        if(XCOUNT == 0x000)
        {
            ledout <= 1;
        }
        if(XCOUNT == ZCOUNT)
        {
            ledout <= 0;
        }


        if(state == 0)
        {
            if(XCOUNT == 0x000)
            {
                ZCOUNT <= ZCOUNT + 1;
            }
            if(ZCOUNT == 0xFFF)
            {
                state <= 1;
            }
        }
        else
        {
            if(XCOUNT == 0x000)
            {
                ZCOUNT <= ZCOUNT - 1;
            }
            if(ZCOUNT == 0x010)
            {
                state <= 0;
            }
        }
        
        LED0 = ledout;
        LED1 = ledout;
        LED2 = ledout;
        LED3 = ledout;
        LED4 = ~ledout;
        LED5 = ~ledout;
        LED6 = ~ledout;
        LED7 = ~ledout;
    }
}
